module B
  (
   input  inA,
   input  inB,
   output outC
   );

assign outC = inA + inB;

endmodule // B
